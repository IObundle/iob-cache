   //General Interface Signals (do not remove indentation)
   //START_IO_TABLE gen
   `IOB_INPUT(clk,          1), //System clock
   `IOB_INPUT(reset,        1), //System reset, asynchronous and active high
