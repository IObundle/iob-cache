//DERIVED MACROS
`define IOB_CACHE_NBYTES (DATA_W/8)
`define IOB_CACHE_NBYTES_W ($clog2(`IOB_CACHE_NBYTES))
`define IOB_CACHE_BE_NBYTES (BE_DATA_W/8)
`define IOB_CACHE_BE_NBYTES_W ($clog2(`IOB_CACHE_BE_NBYTES))
`define IOB_CACHE_LINE2BE_W (WORD_OFFSET_W-$clog2(BE_DATA_W/DATA_W))
