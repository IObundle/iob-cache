//DERIVED MACROS
`define IOB_CACHE_NBYTES (`IOB_CACHE_DATA_W/8)
`define IOB_CACHE_NBYTES_W ($clog2(`IOB_CACHE_NBYTES))
`define IOB_CACHE_BE_NBYTES (`IOB_CACHE_BE_DATA_W/8)
`define IOB_CACHE_BE_NBYTES_W ($clog2(`IOB_CACHE_BE_NBYTES))
`define IOB_CACHE_LINE2BE_W (`IOB_CACHE_WORD_OFFSET_W-$clog2(`IOB_CACHE_BE_DATA_W/`IOB_CACHE_DATA_W))
