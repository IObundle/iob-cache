// SPDX-FileCopyrightText: 2025 IObundle
//
// SPDX-License-Identifier: MIT

`include "iob_uut_conf.vh"
`define IOB_CSRS_ADDR_W (`IOB_UUT_FE_ADDR_W)
