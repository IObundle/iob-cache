`timescale 1ns / 1ps

`include "iob_cache_conf.vh"

module iob_cache_back_end #(
   parameter ADDR_W     = `IOB_CACHE_ADDR_W,
   parameter DATA_W     = `IOB_CACHE_DATA_W,
   parameter BE_ADDR_W     = `IOB_CACHE_BE_ADDR_W,
   parameter BE_DATA_W     = `IOB_CACHE_BE_DATA_W,
   parameter WORD_OFFSET_W = `IOB_CACHE_WORD_OFFSET_W,
   parameter WRITE_POL     = `IOB_CACHE_WRITE_THROUGH,
   parameter WTBUF_DEPTH_W = `IOB_CACHE_WTBUF_DEPTH_W,

   //derived parameters
   parameter FE_NBYTES     = DATA_W / 8,
   parameter FE_NBYTES_W   = $clog2(FE_NBYTES),
   parameter BE_NBYTES     = BE_DATA_W / 8,
   parameter BE_NBYTES_W   = $clog2(BE_NBYTES),
   parameter LINE2BE_W     = WORD_OFFSET_W - $clog2(BE_DATA_W / DATA_W)
) (
   // write channel
   input                                                                        write_req_i,
   input [ ADDR_W-1 : FE_NBYTES_W + WRITE_POL*WORD_OFFSET_W]                 write_addr_i,
   input [DATA_W + WRITE_POL*(DATA_W*(2**WORD_OFFSET_W)-DATA_W)-1 : 0] write_wdata_i,
   input [ FE_NBYTES-1:0]                                                       write_wstrb_i,
   output                                                                       write_ack_o,

   // read channel
   input                                                                        read_req_i,
   input [ADDR_W-1:BE_NBYTES_W + LINE2BE_W]                                  read_addr_i,
   output                                                                       read_valid_o,
   output [ LINE2BE_W -1:0]                                                     read_addr_o,
   output                                                                       read_busy_o,

   // back-end memory interface
   output [ 1-1:0]                                                              be_iob_avalid_o,
   output [ BE_ADDR_W-1:0]                                                      be_iob_addr_o,
   output [ BE_DATA_W-1:0]                                                      be_iob_wdata_o,
   output [(BE_DATA_W/8)-1:0]                                                   be_iob_wstrb_o,
   input [ 1-1:0]                                                               be_iob_rvalid_i,
   input [ BE_DATA_W-1:0]                                                       be_iob_rdata_i,
   input [ 1-1:0]                                                               be_iob_ready_i,
                                                                                
                                                                                `include "iob_clkrst_port.vs"
   );

   wire be_valid_read, be_valid_write;
   assign be_iob_avalid_o = be_valid_read | be_valid_write;

   wire [BE_ADDR_W-1:0] be_addr_read, be_addr_write;
   assign be_iob_addr_o  = (be_valid_read) ? be_addr_read : be_addr_write;

   iob_cache_read_channel #(
      .ADDR_W    (ADDR_W),
      .DATA_W    (DATA_W),
      .BE_ADDR_W    (BE_ADDR_W),
      .BE_DATA_W    (BE_DATA_W),
      .WORD_OFFSET_W(WORD_OFFSET_W)
   ) read_fsm (
      .clk_i       (clk_i),
      .arst_i      (arst_i),
               
      .read_req_i(read_req_i),
      .read_req_addr_i (read_addr_i),
      .read_valid_o(read_valid_o),
      .read_addr_o (read_addr_o),
      .read_busy_o (read_busy_o),

      .be_addr_o   (be_addr_read),
      .be_valid_o  (be_valid_read),
      .be_rvalid_i (be_iob_rvalid_i),
      .be_rdata_i  (be_iob_rdata_i),
      .be_ready_i  (be_iob_ready_i)
   );

   iob_cache_write_channel #(
      .ADDR_W       (ADDR_W),
      .DATA_W       (DATA_W),
      .BE_ADDR_W    (BE_ADDR_W),
      .BE_DATA_W    (BE_DATA_W),
      .WRITE_POL    (WRITE_POL),
      .WORD_OFFSET_W(WORD_OFFSET_W)
   ) write_fsm (
      .clk_i(clk_i),
      .arst_i(arst_i),

      .valid_i(write_req_i),
      .addr_i (write_addr_i),
      .wstrb_i(write_wstrb_i),
      .wdata_i(write_wdata_i),
      .wack_o(write_ack_o),

      .be_valid_o(be_valid_write),
      .be_addr_o (be_addr_write),
      .be_wdata_o(be_iob_wdata_o),
      .be_wstrb_o(be_iob_wstrb_o),
      .be_ready_i(be_iob_ready_i)
   );





   
endmodule
